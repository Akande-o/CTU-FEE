library verilog;
use verilog.vl_types.all;
entity BeaconAEs_vlg_check_tst is
    port(
        M               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end BeaconAEs_vlg_check_tst;
