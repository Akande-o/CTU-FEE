library verilog;
use verilog.vl_types.all;
entity BeaconAE_vlg_vec_tst is
end BeaconAE_vlg_vec_tst;
