library verilog;
use verilog.vl_types.all;
entity BeaconAEs_vlg_vec_tst is
end BeaconAEs_vlg_vec_tst;
